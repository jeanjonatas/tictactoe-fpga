module cpu(matriz , clock);

input matrix;
